
module shifter(
input clk,rst,flag,
output reg [3:0]out
);

//write your code..



endmodule